module controllers

pub struct WebSocket{}
