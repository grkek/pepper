module controllers

pub struct Http {}
